module regm_tb;

    

    Mreg M()

endmodule